-- Generate next state based on curent state and inputs

library STD;
library IEEE;
use IEEE.std_logic_1164.all;

entity next_state_gen is

end next_state_gen;

architecture structural of next_state_gen is

begin

end structural;

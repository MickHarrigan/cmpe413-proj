library STD;
library IEEE;
use IEEE.std_logic_1164.all;

entity encoder32to5 is
    port(
        input0      : in std_logic;
        input1      : in std_logic;
        input2      : in std_logic;
        input3      : in std_logic;
        input4      : in std_logic;
        input5      : in std_logic;
        input6      : in std_logic;
        input7      : in std_logic;
        input8      : in std_logic;
        input9      : in std_logic;
        input10     : in std_logic;
        input11     : in std_logic;
        input12     : in std_logic;
        input13     : in std_logic;
        input14     : in std_logic;
        input15     : in std_logic;
        input16     : in std_logic;
        input17     : in std_logic;
        input18     : in std_logic;
        input19     : in std_logic;
        input20     : in std_logic;
        input21     : in std_logic;
        input22     : in std_logic;
        input23     : in std_logic;
        input24     : in std_logic;
        input25     : in std_logic;
        input26     : in std_logic;
        input27     : in std_logic;
        input28     : in std_logic;
        input29     : in std_logic;
        input30     : in std_logic;
        input31     : in std_logic;
        output0     : out std_logic_vector(4 downto 0);
    );
end encoder32to5;